../../../TheSDK_generators/verilog/f2_dsp.v