../../../TheSDK_generators/verilog/tb_f2_dsp.v