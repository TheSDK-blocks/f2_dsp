../chisel/verilog/f2_dsp.v