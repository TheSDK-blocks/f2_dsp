../../../TheSDK_generators/f2_dsp_and_serdes/f2_dsp/verilog/f2_dsp.v